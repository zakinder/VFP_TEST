package frame_en_lib;
    `define sbmsbl_v1                      1
endpackage
