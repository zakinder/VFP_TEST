package frame_en_lib;
    `define rgb_v1                      1
endpackage
