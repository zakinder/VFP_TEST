package frame_en_lib;
    `define emboss_v3                      1
endpackage
