package frame_en_lib;
    `define hsv_v0                      1
endpackage
