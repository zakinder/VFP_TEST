package frame_en_lib;
    `define sharp_v2                      1
endpackage
