package frame_en_lib;
    `define cgain_v0                      1
endpackage
