package frame_en_lib;
    `define cgain_v3                      1
endpackage
