// MODULE : VFPCONFIGDUT
module vfpConfigDut(axi4l_if.ConfigMaster axi4l_vif,axi4s_if.rx_channel axi4s_vif,tp_if.templateSlave tp_vif,d5m_camera_if.ConfigMaster d5m_camera_vif);
import generic_pack::*;  
    VFP_v1_0                  #(
    .revision_number           ( revision_number            ),
    .C_rgb_m_axis_TDATA_WIDTH  ( C_rgb_m_axis_TDATA_WIDTH   ),
    .C_rgb_m_axis_START_COUNT  ( C_rgb_m_axis_START_COUNT   ),
    .C_rgb_s_axis_TDATA_WIDTH  ( C_rgb_s_axis_TDATA_WIDTH   ),
    .C_m_axis_mm2s_TDATA_WIDTH ( C_m_axis_mm2s_TDATA_WIDTH  ),
    .C_m_axis_mm2s_START_COUNT ( C_m_axis_mm2s_START_COUNT  ),
    .C_vfpConfig_DATA_WIDTH    ( C_vfpConfig_DATA_WIDTH     ),
    .C_vfpConfig_ADDR_WIDTH    ( C_vfpConfig_ADDR_WIDTH     ),
    .conf_data_width           ( conf_data_width            ),
    .conf_addr_width           ( conf_addr_width            ),
    .i_data_width              ( i_data_width               ),
    .s_data_width              ( s_data_width               ),
    .b_data_width              ( b_data_width               ),
    .i_precision               ( i_precision                ),
    .i_full_range              ( i_full_range               ),
    .img_width                 ( img_width                  ),
    .dataWidth                 ( dataWidth                  ))
    dutVFP_v1Inst              (
    //d5m input
    .pixclk                    (d5m_camera_vif.pixclk        ),//(d5m_camera_vif.ACLK   ),
    .ifval                     (d5m_camera_vif.ifval         ),//(d5m_camera_vif.ARESETN),
    .ilval                     (d5m_camera_vif.ilval         ),//(d5m_camera_vif.AWADDR ),
    .idata                     (d5m_camera_vif.idata         ),//(d5m_camera_vif.AWPROT ),
    //tx channel
    .rgb_m_axis_aclk           (axi4s_vif.ACLK               ),
    .rgb_m_axis_aresetn        (axi4s_vif.ARESET_N           ),
    .rgb_m_axis_tready         (                             ),//(axi4l_vif.AWADDR ),
    .rgb_m_axis_tvalid         (                             ),//(axi4l_vif.AWPROT ),
    .rgb_m_axis_tlast          (                             ),//(axi4l_vif.AWVALID),
    .rgb_m_axis_tuser          (                             ),//(axi4l_vif.AWREADY),
    .rgb_m_axis_tdata          (                             ),//(axi4l_vif.WDATA  ),
    //rx channel               
    .rgb_s_axis_aclk           (axi4s_vif.ACLK               ),
    .rgb_s_axis_aresetn        (axi4s_vif.ARESET_N           ),
    .rgb_s_axis_tready         (axi4s_vif.TREADY             ),
    .rgb_s_axis_tvalid         (axi4s_vif.TVALID             ),
    .rgb_s_axis_tlast          (axi4s_vif.TLAST              ),
    .rgb_s_axis_tuser          (axi4s_vif.TUSER              ),
    .rgb_s_axis_tdata          (axi4s_vif.TDATA              ),
    //destination channel                                    
    .m_axis_mm2s_aclk          (axi4s_vif.ACLK               ),
    .m_axis_mm2s_aresetn       (axi4s_vif.ARESET_N           ),
    .m_axis_mm2s_tready        (                             ),//(axi4l_vif.AWADDR ),
    .m_axis_mm2s_tvalid        (                             ),//(axi4l_vif.AWPROT ),
    .m_axis_mm2s_tuser         (                             ),//(axi4l_vif.AWVALID),
    .m_axis_mm2s_tlast         (                             ),//(axi4l_vif.AWREADY),
    .m_axis_mm2s_tdata         (                             ),//(axi4l_vif.WDATA  ),
    .m_axis_mm2s_tkeep         (                             ),//(axi4l_vif.AWPROT ),
    .m_axis_mm2s_tstrb         (                             ),//(axi4l_vif.AWVALID),
    .m_axis_mm2s_tid           (                             ),//(axi4l_vif.AWREADY),
    .m_axis_mm2s_tdest         (                             ),//(axi4l_vif.WDATA  ),
    //video configuration      
    .vfpconfig_aclk            (axi4l_vif.ACLK               ),
    .vfpconfig_aresetn         (axi4l_vif.ARESETN            ),
    .vfpconfig_awaddr          (axi4l_vif.AWADDR             ),
    .vfpconfig_awprot          (axi4l_vif.AWPROT             ),
    .vfpconfig_awvalid         (axi4l_vif.AWVALID            ),
    .vfpconfig_awready         (axi4l_vif.AWREADY            ),
    .vfpconfig_wdata           (axi4l_vif.WDATA              ),
    .vfpconfig_wstrb           (axi4l_vif.WSTRB              ),
    .vfpconfig_wvalid          (axi4l_vif.WVALID             ),
    .vfpconfig_wready          (axi4l_vif.WREADY             ),
    .vfpconfig_bresp           (axi4l_vif.BRESP              ),
    .vfpconfig_bvalid          (axi4l_vif.BVALID             ),
    .vfpconfig_bready          (axi4l_vif.BREADY             ),
    .vfpconfig_araddr          (axi4l_vif.ARADDR             ),
    .vfpconfig_arprot          (axi4l_vif.ARPROT             ),
    .vfpconfig_arvalid         (axi4l_vif.ARVALID            ),
    .vfpconfig_arready         (axi4l_vif.ARREADY            ),
    .vfpconfig_rdata           (axi4l_vif.RDATA              ),
    .vfpconfig_rresp           (axi4l_vif.RRESP              ),
    .vfpconfig_rvalid          (axi4l_vif.RVALID             ),
    .vfpconfig_rready          (axi4l_vif.RREADY             ));
endmodule: vfpConfigDut