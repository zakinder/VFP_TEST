package frame_en_lib;
    `define sharp_v0                      1
endpackage
