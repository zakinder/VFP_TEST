package frame_en_lib;
    `define sobel_v0                      1
endpackage
