package frame_en_lib;
    `define rgb_v0                      1
endpackage
