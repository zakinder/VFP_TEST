package frame_en_lib;
    `define hsl_v0                      1
endpackage
