package frame_en_lib;
    `define hsv_v2                      1
endpackage
