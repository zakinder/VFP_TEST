package frame_en_lib;
    `define sbmsbl_v0                      1
endpackage
