package frame_en_lib;
    `define cgtocg_v1                      1
endpackage
