package frame_en_lib;
    `define emboss_v0    1
endpackage
