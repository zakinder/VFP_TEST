// Class: d5m_camera_configuration
class d5m_camera_configuration extends uvm_object;
    `uvm_object_utils(d5m_camera_configuration)
    // Function: new
    function new(string name = "");
        super.new(name);
    endfunction: new
endclass: d5m_camera_configuration