  `include "../../agents/d5m_agent/d5m_camera_agent_pkg.sv"
package d5m_camera_pkg;
  import d5m_camera_agent_pkg::*;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  `include "../../defin_lib.svh"
  `include "d5m_camera_env.sv"
  `include "../../test/d5m_camera/d5m_camera_test.sv"
  `include "../../test/d5m_camera/d5m_camera_image_pattern_test.sv"
  `include "../../test/d5m_camera/d5m_camera_image_file_test.sv"
  `include "../../test/d5m_camera/d5m_rgb_patten_test.sv"
endpackage:d5m_camera_pkg
