    `define cgtocg_v1                      1
endpackage
