package frame_en_lib;
    `define cgain_v2                      1
endpackage
