package frame_en_lib;
    `define sobel_v2                      1
endpackage
