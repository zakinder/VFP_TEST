package frame_en_lib;
    `define sbmshl_v0                      1
endpackage
