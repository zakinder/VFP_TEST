package frame_en_lib;
    `define sbmshl_v1                      1
endpackage
